module beat32 (


);

endmodule