module master_fsm_tb ();


endmodule