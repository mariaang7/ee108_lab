module sine_reader (
// TODO: fill in your implementation from lab 4! 

);

endmodule