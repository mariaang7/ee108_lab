module verifier
