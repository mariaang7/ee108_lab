module float_add_tb (

);

// your implementation goes here!



endmodule