module big_number_first (

);

// your implementation goes here!



endmodule