module bicycle_fsm_tb ();


endmodule