module shifter (

);

// your implementation goes here!



endmodule