module master_fsm (

);


endmodule