module beat32_tb ();


endmodule