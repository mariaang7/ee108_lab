module blinker (

);


endmodule