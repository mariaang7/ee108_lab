module shifter (

);

endmodule