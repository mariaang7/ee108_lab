module programmable_blinker (
  Input wire shift_left, shift_right,
  output wire out
);

  shifter jeff (.shift_left(shift_left), .shift_right(shift_right), 
 

endmodule
