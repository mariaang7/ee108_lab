module hasher (
  input wire [63:0] username,
  input wire [63:0] password,
  output wire valid
);
