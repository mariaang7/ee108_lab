module song_rom (
// TODO: fill in your implementation from lab 4! 

);

endmodule