module timer (

);


endmodule