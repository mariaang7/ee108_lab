module adder_tb (

);

// your implementation goes here!



endmodule