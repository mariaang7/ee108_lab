module programmable_blinker (

);


endmodule