module master_fsm (input 

);


endmodule
