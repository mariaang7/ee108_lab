module shifter_tb ();

endmodule