module mcu (
// TODO: fill in your implementation from lab 4! 

);

endmodule