module big_number_first_tb (

);

// your implementation goes here!



endmodule