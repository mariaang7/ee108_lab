module shifter_tb (

);

// your implementation goes here!



endmodule