module adder (

);

// your implementation goes here!



endmodule