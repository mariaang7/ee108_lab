module programmable_blinker_tb ();

endmodule