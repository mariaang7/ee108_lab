module master_fsm (input wire next;
                   input wire slower;
                   input wire faster;

);


endmodule
