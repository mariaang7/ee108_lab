module blinker_tb ();

endmodule