module hasher
