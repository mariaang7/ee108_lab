module timer_tb ();

endmodule 